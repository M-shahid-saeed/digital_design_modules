interface multiplier_intf #(parameter N=8) (input logic clk);
  logic [N-1:0] Data_in_A;
  logic [N-1:0] Data_in_B;
  logic Reset;      
  logic EA, EB;     
  logic [(2*N)-1:0] P_out; 
endinterface